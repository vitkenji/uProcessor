library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ROM is
port(
    clk : in std_logic;
    address : in unsigned(6 downto 0);
    data : out unsigned(16 downto 0)
);
end entity;

architecture ROM_arch of ROM is
    type mem is array (0 to 127) of unsigned(16 downto 0);
    constant ROM_content : mem := (
        0   => "00000000000000000",
        1   => "00000000000000001",
        2   => "00000000000000010",
        3   => "00000000000000011",
        4   => "00000000000000100",
        5   => "00000000000000101",
        6   => "00000000000000110",
        7   => "00000000000000111",
        8   => "00000000000001000",
        9   => "00000000000001001",
        10  => "00000000000001010",
        11  => "00000000000001011",
        12  => "00000000000001100",
        13  => "00000000000001101",
        14  => "00000000000001110",
        15  => "00000000000001111",
        16  => "00000000000010000",
        17  => "00000000000010001",
        18  => "00000000000010010",
        19  => "00000000000010011",
        20  => "00000000000010100",
        21  => "00000000000010101",
        22  => "00000000000010110",
        23  => "00000000000010111",
        24  => "00000000000011000",
        25  => "00000000000011001",
        26  => "00000000000011010",
        27  => "00000000000011011",
        28  => "00000000000011100",
        29  => "00000000000011101",
        30  => "00000000000011110",
        31  => "00000000000011111",
        32  => "00000000000100000",
        33  => "00000000000100001",
        34  => "00000000000100010",
        35  => "00000000000100011",
        36  => "00000000000100100",
        37  => "00000000000100101",
        38  => "00000000000100110",
        39  => "00000000000100111",
        40  => "00000000000101000",
        others => (others =>'0')
    );
    begin
        process(clk)
        begin
            if (rising_edge(clk)) then
                data <= ROM_content(to_integer(address));
            end if;
        end process;
end architecture;