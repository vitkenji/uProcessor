library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity State_Machine_tb is
end;

architecture State_Machine_tb_arch of State_Machine_tb is
    process
    begin
    end process;
end architecture;

