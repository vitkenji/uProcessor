library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity Control_Unit is
    port(

    );
end entity;

architecture Control_Unit_arch of Control_Unit is
end architecture;