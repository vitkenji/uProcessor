library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity PC is
    port (

    );
end entity;

architecture PC_arch of PC is
end architecture;