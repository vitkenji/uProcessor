library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity State_Machine is
    port(

    );
end entity;

architecture State_Machine_arch of State_Machine is
    process
    begin
    end process;
end architecture;