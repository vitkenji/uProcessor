library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity Control_Unit_tb is
end;

architecture Control_Unit_tb_arch of Control_Unit_tb is
    
end architecture;