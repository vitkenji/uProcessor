library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- Operações da ALU
-- 00 -> soma [1+0 = 1; 0+1 = 1; 0+0 = 0; 1+1 = 10;]
-- 01 -> subtração [1-0 = 1; 0-1 = 1; 1-1 = 0; 0-0 = 0]
-- 10 -> and [Aplica a operação and bit a bit entre os dois números]
-- 11 -> xor [Aplica a operação xor bit a bit entre os dois números]

entity ALU is
    port (
        input_0, input_1 : in unsigned (15 downto 0);
        operation_selector: in unsigned (1 downto 0);
        carry, greater_equal, less_equal: out std_logic; 
        saida : out unsigned (15 downto 0)
    );
end entity;

architecture ALU_arch of ALU is

    -- Sinais auxiliares
    signal input_0_17bits, input_1_17bits, sum_result, sub_result : unsigned(16 downto 0);

begin
    -- [*] Melhoria Futura: Tratamento com números negativos, ou seja, não usar mais unsigned e sim como signed
    input_0 <= unsigned(input_0);
    input_1 <= unsigned(input_1);

    -- Formando 17 bits para armazenar o carry junto com o resultado da operação
    input_0_17bits <= '0' & input_0;
    input_1_17bits <= '0' & input_1;

    sum_result_17bits <= input_0_17bits + input_1_17bits; -- Carry
    sub_result_17bits <= input_0_17bits - input_1_17bits; -- Borrow

    saida <= input_0 + input_1 when operation_selector = "00" else
              input_0 - input_1 when operation_selector = "01" else
              input_0 and input_1 when operation_selector = "10" else
              input_0 xor input_1 when operation_selector = "11" else
              "0000000000000000";

    carry <= sum_result_17bits(16) when operation_selector = "00" else
             sub_result_17bits(16) when operation_selector = "01" else
             '0';

    greater_equal <= '1' when input_0 >= input_1 else '0';
    less_equal <= '1' when input_0 <= input_1 else '0';

end architecture;